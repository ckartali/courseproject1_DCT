`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 14.04.2024 11:38:55
// Design Name: 
// Module Name: tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module tb();

reg [14:0] in;
wire [17:0] out1,out2,out3,out4;
reg clk;
reg rst;


add_up x2(in,out1,out2,out4,out3,clk,rst);

initial clk=1'b1;
always #1 clk=~clk;

initial
begin
rst=1'b1;

#20
rst=1'b0;
//in=13'b000_1000000000;
//#2 in=13'b000_1000000000;
//#2 in=13'b000_1000000000;
//#2 in=13'b000_1000000000;
//#2 in=13'b000_1000000000;
//#2 in=13'b000_1000000000;
//#2 in=13'b000_1000000000;
//#2 in=13'b000_1000000000;
//#2 in=13'b000_1000000000;
//#2 in=13'b000_1000000000;
//#2 in=13'b000_1000000000;
//#2 in=13'b000_1000000000;
//#2 in=13'b000_1000000000;
//#2 in=13'b000_1000000000;
//#2 in=13'b000_1000000000;
//#2 in=13'b000_1000000000;
//in=13'b111_1000000000;
//#2 in=13'b111_1000000000;
//#2 in=13'b111_1000000000;
//#2 in=13'b111_1000000000;
//#2 in=13'b111_1000000000;
//#2 in=13'b111_1000000000;
//#2 in=13'b111_1000000000;
//#2 in=13'b111_1000000000;
//#2 in=13'b111_1000000000;
//#2 in=13'b111_1000000000;
//#2 in=13'b111_1000000000;
//#2 in=13'b111_1000000000;
//#2 in=13'b111_1000000000;
//#2 in=13'b111_1000000000;
//#2 in=13'b111_1000000000;
//#2 in=13'b111_1000000000;
in=15'b00001_0000000000;
#2 in=15'b00010_0000000000;
#2 in=15'b00011_0000000000;
#2 in=15'b00100_0000000000;
#2 in=15'b00101_0000000000;
#2 in=15'b00110_0000000000;
#2 in=15'b00111_0000000000;
#2 in=15'b01000_0000000000;
#2 in=15'b01001_0000000000;
#2 in=15'b00001_1000000000;
#2 in=15'b00010_1000000000;
#2 in=15'b00011_1000000000;
#2 in=15'b00100_1000000000;
#2 in=15'b00101_1000000000;
#2 in=15'b00110_1000000000;
#2 in=15'b00111_1000000000;



#500 $finish;
end
endmodule
