`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 19.04.2024 21:38:12
// Design Name: 
// Module Name: ROM4
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module ROM4(
   input [7:0] A,input [2:0]k,

    output reg [14:0] out
    );

//storing for X3,X7,X11,X15    
always @ (*)
begin
    if (k==0) 
        begin
            if(A==8'd0)
                out<=15'b000000000000000;
            else if(A==8'd1)
                out<=15'b111111011010111;
            else if(A==8'd2)
                out<=15'b111110011101001;
            else if(A==8'd3)
                out<=15'b111101111000000;
            else if(A==8'd4)
                out<=15'b111110000000101;
            else if(A==8'd5)
                out<=15'b111101011011100;
            else if(A==8'd6)
                out<=15'b111100011101110;
            else if(A==8'd7)
                out<=15'b111011111000101;
            else if(A==8'd8)
                out<=15'b111110001111001;
            else if(A==8'd9)
                out<=15'b111101101010000;
            else if(A==8'd10)
                out<=15'b111100101100010;
            else if(A==8'd11)
                out<=15'b111100000111001;
            else if(A==8'd12)
                out<=15'b111100001111110;
            else if(A==8'd13)
                out<=15'b111011101010101;
            else if(A==8'd14)
                out<=15'b111010101100111;
            else if(A==8'd15)
                out<=15'b111010000111110;
            else if(A==8'd16)
                out<=15'b111111000011110;
            else if(A==8'd17)
                out<=15'b111110011110101;
            else if(A==8'd18)
                out<=15'b111101100000111;
            else if(A==8'd19)
                out<=15'b111100111011110;
            else if(A==8'd20)
                out<=15'b111101000100011;
            else if(A==8'd21)
                out<=15'b111100011111010;
            else if(A==8'd22)
                out<=15'b111011100001100;
            else if(A==8'd23)
                out<=15'b111010111100011;
            else if(A==8'd24)
                out<=15'b111101010010111;
            else if(A==8'd25)
                out<=15'b111100101101110;
            else if(A==8'd26)
                out<=15'b111011110000000;
            else if(A==8'd27)
                out<=15'b111011001010111;
            else if(A==8'd28)
                out<=15'b111011010011100;
            else if(A==8'd29)
                out<=15'b111010101110011;
            else if(A==8'd30)
                out<=15'b111001110000101;
            else if(A==8'd31)
                out<=15'b111001001011100;
            else if(A==8'd32)
                out<=15'b000000001100100;
            else if(A==8'd33)
                out<=15'b111111100111011;
            else if(A==8'd34)
                out<=15'b111110101001101;
            else if(A==8'd35)
                out<=15'b111110000100100;
            else if(A==8'd36)
                out<=15'b111110001101001;
            else if(A==8'd37)
                out<=15'b111101101000000;
            else if(A==8'd38)
                out<=15'b111100101010010;
            else if(A==8'd39)
                out<=15'b111100000101001;
            else if(A==8'd40)
                out<=15'b111110011011101;
            else if(A==8'd41)
                out<=15'b111101110110100;
            else if(A==8'd42)
                out<=15'b111100111000110;
            else if(A==8'd43)
                out<=15'b111100010011101;
            else if(A==8'd44)
                out<=15'b111100011100010;
            else if(A==8'd45)
                out<=15'b111011110111001;
            else if(A==8'd46)
                out<=15'b111010111001011;
            else if(A==8'd47)
                out<=15'b111010010100010;
            else if(A==8'd48)
                out<=15'b111111010000010;
            else if(A==8'd49)
                out<=15'b111110101011001;
            else if(A==8'd50)
                out<=15'b111101101101011;
            else if(A==8'd51)
                out<=15'b111101001000010;
            else if(A==8'd52)
                out<=15'b111101010000111;
            else if(A==8'd53)
                out<=15'b111100101011110;
            else if(A==8'd54)
                out<=15'b111011101110000;
            else if(A==8'd55)
                out<=15'b111011001000111;
            else if(A==8'd56)
                out<=15'b111101011111011;
            else if(A==8'd57)
                out<=15'b111100111010010;
            else if(A==8'd58)
                out<=15'b111011111100100;
            else if(A==8'd59)
                out<=15'b111011010111011;
            else if(A==8'd60)
                out<=15'b111011100000000;
            else if(A==8'd61)
                out<=15'b111010111010111;
            else if(A==8'd62)
                out<=15'b111001111101001;
            else if(A==8'd63)
                out<=15'b111001011000000;
            else if(A==8'd64)
                out<=15'b000001010001001;
            else if(A==8'd65)
                out<=15'b000000101100000;
            else if(A==8'd66)
                out<=15'b111111101110010;
            else if(A==8'd67)
                out<=15'b111111001001001;
            else if(A==8'd68)
                out<=15'b111111010001110;
            else if(A==8'd69)
                out<=15'b111110101100101;
            else if(A==8'd70)
                out<=15'b111101101110111;
            else if(A==8'd71)
                out<=15'b111101001001110;
            else if(A==8'd72)
                out<=15'b111111100000010;
            else if(A==8'd73)
                out<=15'b111110111011001;
            else if(A==8'd74)
                out<=15'b111101111101011;
            else if(A==8'd75)
                out<=15'b111101011000010;
            else if(A==8'd76)
                out<=15'b111101100000111;
            else if(A==8'd77)
                out<=15'b111100111011110;
            else if(A==8'd78)
                out<=15'b111011111110000;
            else if(A==8'd79)
                out<=15'b111011011000111;
            else if(A==8'd80)
                out<=15'b000000010100111;
            else if(A==8'd81)
                out<=15'b111111101111110;
            else if(A==8'd82)
                out<=15'b111110110010000;
            else if(A==8'd83)
                out<=15'b111110001100111;
            else if(A==8'd84)
                out<=15'b111110010101100;
            else if(A==8'd85)
                out<=15'b111101110000011;
            else if(A==8'd86)
                out<=15'b111100110010101;
            else if(A==8'd87)
                out<=15'b111100001101100;
            else if(A==8'd88)
                out<=15'b111110100100000;
            else if(A==8'd89)
                out<=15'b111101111110111;
            else if(A==8'd90)
                out<=15'b111101000001001;
            else if(A==8'd91)
                out<=15'b111100011100000;
            else if(A==8'd92)
                out<=15'b111100100100101;
            else if(A==8'd93)
                out<=15'b111011111111100;
            else if(A==8'd94)
                out<=15'b111011000001110;
            else if(A==8'd95)
                out<=15'b111010011100101;
            else if(A==8'd96)
                out<=15'b000001011101101;
            else if(A==8'd97)
                out<=15'b000000111000100;
            else if(A==8'd98)
                out<=15'b111111111010110;
            else if(A==8'd99)
                out<=15'b111111010101101;
            else if(A==8'd100)
                out<=15'b111111011110010;
            else if(A==8'd101)
                out<=15'b111110111001001;
            else if(A==8'd102)
                out<=15'b111101111011011;
            else if(A==8'd103)
                out<=15'b111101010110010;
            else if(A==8'd104)
                out<=15'b111111101100110;
            else if(A==8'd105)
                out<=15'b111111000111101;
            else if(A==8'd106)
                out<=15'b111110001001111;
            else if(A==8'd107)
                out<=15'b111101100100110;
            else if(A==8'd108)
                out<=15'b111101101101011;
            else if(A==8'd109)
                out<=15'b111101001000010;
            else if(A==8'd110)
                out<=15'b111100001010100;
            else if(A==8'd111)
                out<=15'b111011100101011;
            else if(A==8'd112)
                out<=15'b000000100001011;
            else if(A==8'd113)
                out<=15'b111111111100010;
            else if(A==8'd114)
                out<=15'b111110111110100;
            else if(A==8'd115)
                out<=15'b111110011001011;
            else if(A==8'd116)
                out<=15'b111110100010000;
            else if(A==8'd117)
                out<=15'b111101111100111;
            else if(A==8'd118)
                out<=15'b111100111111001;
            else if(A==8'd119)
                out<=15'b111100011010000;
            else if(A==8'd120)
                out<=15'b111110110000100;
            else if(A==8'd121)
                out<=15'b111110001011011;
            else if(A==8'd122)
                out<=15'b111101001101101;
            else if(A==8'd123)
                out<=15'b111100101000100;
            else if(A==8'd124)
                out<=15'b111100110001001;
            else if(A==8'd125)
                out<=15'b111100001100000;
            else if(A==8'd126)
                out<=15'b111011001110010;
            else if(A==8'd127)
                out<=15'b111010101001001;
            else if(A==8'd128)
                out<=15'b000001111010011;
            else if(A==8'd129)
                out<=15'b000001010101010;
            else if(A==8'd130)
                out<=15'b000000010111100;
            else if(A==8'd131)
                out<=15'b111111110010011;
            else if(A==8'd132)
                out<=15'b111111111011000;
            else if(A==8'd133)
                out<=15'b111111010101111;
            else if(A==8'd134)
                out<=15'b111110011000001;
            else if(A==8'd135)
                out<=15'b111101110011000;
            else if(A==8'd136)
                out<=15'b000000001001100;
            else if(A==8'd137)
                out<=15'b111111100100011;
            else if(A==8'd138)
                out<=15'b111110100110101;
            else if(A==8'd139)
                out<=15'b111110000001100;
            else if(A==8'd140)
                out<=15'b111110001010001;
            else if(A==8'd141)
                out<=15'b111101100101000;
            else if(A==8'd142)
                out<=15'b111100100111010;
            else if(A==8'd143)
                out<=15'b111100000010001;
            else if(A==8'd144)
                out<=15'b000000111110001;
            else if(A==8'd145)
                out<=15'b000000011001000;
            else if(A==8'd146)
                out<=15'b111111011011010;
            else if(A==8'd147)
                out<=15'b111110110110001;
            else if(A==8'd148)
                out<=15'b111110111110110;
            else if(A==8'd149)
                out<=15'b111110011001101;
            else if(A==8'd150)
                out<=15'b111101011011111;
            else if(A==8'd151)
                out<=15'b111100110110110;
            else if(A==8'd152)
                out<=15'b111111001101010;
            else if(A==8'd153)
                out<=15'b111110101000001;
            else if(A==8'd154)
                out<=15'b111101101010011;
            else if(A==8'd155)
                out<=15'b111101000101010;
            else if(A==8'd156)
                out<=15'b111101001101111;
            else if(A==8'd157)
                out<=15'b111100101000110;
            else if(A==8'd158)
                out<=15'b111011101011000;
            else if(A==8'd159)
                out<=15'b111011000101111;
            else if(A==8'd160)
                out<=15'b000010000110111;
            else if(A==8'd161)
                out<=15'b000001100001110;
            else if(A==8'd162)
                out<=15'b000000100100000;
            else if(A==8'd163)
                out<=15'b111111111110111;
            else if(A==8'd164)
                out<=15'b000000000111100;
            else if(A==8'd165)
                out<=15'b111111100010011;
            else if(A==8'd166)
                out<=15'b111110100100101;
            else if(A==8'd167)
                out<=15'b111101111111100;
            else if(A==8'd168)
                out<=15'b000000010110000;
            else if(A==8'd169)
                out<=15'b111111110000111;
            else if(A==8'd170)
                out<=15'b111110110011001;
            else if(A==8'd171)
                out<=15'b111110001110000;
            else if(A==8'd172)
                out<=15'b111110010110101;
            else if(A==8'd173)
                out<=15'b111101110001100;
            else if(A==8'd174)
                out<=15'b111100110011110;
            else if(A==8'd175)
                out<=15'b111100001110101;
            else if(A==8'd176)
                out<=15'b000001001010101;
            else if(A==8'd177)
                out<=15'b000000100101100;
            else if(A==8'd178)
                out<=15'b111111100111110;
            else if(A==8'd179)
                out<=15'b111111000010101;
            else if(A==8'd180)
                out<=15'b111111001011010;
            else if(A==8'd181)
                out<=15'b111110100110001;
            else if(A==8'd182)
                out<=15'b111101101000011;
            else if(A==8'd183)
                out<=15'b111101000011010;
            else if(A==8'd184)
                out<=15'b111111011001110;
            else if(A==8'd185)
                out<=15'b111110110100101;
            else if(A==8'd186)
                out<=15'b111101110110111;
            else if(A==8'd187)
                out<=15'b111101010001110;
            else if(A==8'd188)
                out<=15'b111101011010011;
            else if(A==8'd189)
                out<=15'b111100110101010;
            else if(A==8'd190)
                out<=15'b111011110111100;
            else if(A==8'd191)
                out<=15'b111011010010011;
            else if(A==8'd192)
                out<=15'b000011001011100;
            else if(A==8'd193)
                out<=15'b000010100110011;
            else if(A==8'd194)
                out<=15'b000001101000101;
            else if(A==8'd195)
                out<=15'b000001000011100;
            else if(A==8'd196)
                out<=15'b000001001100001;
            else if(A==8'd197)
                out<=15'b000000100111000;
            else if(A==8'd198)
                out<=15'b111111101001010;
            else if(A==8'd199)
                out<=15'b111111000100001;
            else if(A==8'd200)
                out<=15'b000001011010101;
            else if(A==8'd201)
                out<=15'b000000110101100;
            else if(A==8'd202)
                out<=15'b111111110111110;
            else if(A==8'd203)
                out<=15'b111111010010101;
            else if(A==8'd204)
                out<=15'b111111011011010;
            else if(A==8'd205)
                out<=15'b111110110110001;
            else if(A==8'd206)
                out<=15'b111101111000011;
            else if(A==8'd207)
                out<=15'b111101010011010;
            else if(A==8'd208)
                out<=15'b000010001111010;
            else if(A==8'd209)
                out<=15'b000001101010001;
            else if(A==8'd210)
                out<=15'b000000101100011;
            else if(A==8'd211)
                out<=15'b000000000111010;
            else if(A==8'd212)
                out<=15'b000000001111111;
            else if(A==8'd213)
                out<=15'b111111101010110;
            else if(A==8'd214)
                out<=15'b111110101101000;
            else if(A==8'd215)
                out<=15'b111110000111111;
            else if(A==8'd216)
                out<=15'b000000011110011;
            else if(A==8'd217)
                out<=15'b111111111001010;
            else if(A==8'd218)
                out<=15'b111110111011100;
            else if(A==8'd219)
                out<=15'b111110010110011;
            else if(A==8'd220)
                out<=15'b111110011111000;
            else if(A==8'd221)
                out<=15'b111101111001111;
            else if(A==8'd222)
                out<=15'b111100111100001;
            else if(A==8'd223)
                out<=15'b111100010111000;
            else if(A==8'd224)
                out<=15'b000011011000000;
            else if(A==8'd225)
                out<=15'b000010110010111;
            else if(A==8'd226)
                out<=15'b000001110101001;
            else if(A==8'd227)
                out<=15'b000001010000000;
            else if(A==8'd228)
                out<=15'b000001011000101;
            else if(A==8'd229)
                out<=15'b000000110011100;
            else if(A==8'd230)
                out<=15'b111111110101110;
            else if(A==8'd231)
                out<=15'b111111010000101;
            else if(A==8'd232)
                out<=15'b000001100111001;
            else if(A==8'd233)
                out<=15'b000001000010000;
            else if(A==8'd234)
                out<=15'b000000000100010;
            else if(A==8'd235)
                out<=15'b111111011111001;
            else if(A==8'd236)
                out<=15'b111111100111110;
            else if(A==8'd237)
                out<=15'b111111000010101;
            else if(A==8'd238)
                out<=15'b111110000100111;
            else if(A==8'd239)
                out<=15'b111101011111110;
            else if(A==8'd240)
                out<=15'b000010011011110;
            else if(A==8'd241)
                out<=15'b000001110110101;
            else if(A==8'd242)
                out<=15'b000000111000111;
            else if(A==8'd243)
                out<=15'b000000010011110;
            else if(A==8'd244)
                out<=15'b000000011100011;
            else if(A==8'd245)
                out<=15'b111111110111010;
            else if(A==8'd246)
                out<=15'b111110111001100;
            else if(A==8'd247)
                out<=15'b111110010100011;
            else if(A==8'd248)
                out<=15'b000000101010111;
            else if(A==8'd249)
                out<=15'b000000000101110;
            else if(A==8'd250)
                out<=15'b111111001000000;
            else if(A==8'd251)
                out<=15'b111110100010111;
            else if(A==8'd252)
                out<=15'b111110101011100;
            else if(A==8'd253)
                out<=15'b111110000110011;
            else if(A==8'd254)
                out<=15'b111101001000101;
            else
                out<=15'b111100100011100;
        end 
    
    else if(k==1)
        begin
            if(A==8'd0)
                out<=15'b000000000000000;
            else if(A==8'd1)
                out<=15'b111110101110111;
            else if(A==8'd2)
                out<=15'b111110001111001;
            else if(A==8'd3)
                out<=15'b111100111110000;
            else if(A==8'd4)
                out<=15'b000000100101001;
            else if(A==8'd5)
                out<=15'b111111010100000;
            else if(A==8'd6)
                out<=15'b111110110100010;
            else if(A==8'd7)
                out<=15'b111101100011001;
            else if(A==8'd8)
                out<=15'b000001111111011;
            else if(A==8'd9)
                out<=15'b000000101110010;
            else if(A==8'd10)
                out<=15'b000000001110100;
            else if(A==8'd11)
                out<=15'b111110111101011;
            else if(A==8'd12)
                out<=15'b000010100100100;
            else if(A==8'd13)
                out<=15'b000001010011011;
            else if(A==8'd14)
                out<=15'b000000110011101;
            else if(A==8'd15)
                out<=15'b111111100010100;
            else if(A==8'd16)
                out<=15'b000000001100100;
            else if(A==8'd17)
                out<=15'b111110111011011;
            else if(A==8'd18)
                out<=15'b111110011011101;
            else if(A==8'd19)
                out<=15'b111101001010100;
            else if(A==8'd20)
                out<=15'b000000110001101;
            else if(A==8'd21)
                out<=15'b111111100000100;
            else if(A==8'd22)
                out<=15'b111111000000110;
            else if(A==8'd23)
                out<=15'b111101101111101;
            else if(A==8'd24)
                out<=15'b000010001011111;
            else if(A==8'd25)
                out<=15'b000000111010110;
            else if(A==8'd26)
                out<=15'b000000011011000;
            else if(A==8'd27)
                out<=15'b111111001001111;
            else if(A==8'd28)
                out<=15'b000010110001000;
            else if(A==8'd29)
                out<=15'b000001011111111;
            else if(A==8'd30)
                out<=15'b000001000000001;
            else if(A==8'd31)
                out<=15'b111111101111000;
            else if(A==8'd32)
                out<=15'b111110000101101;
            else if(A==8'd33)
                out<=15'b111100110100100;
            else if(A==8'd34)
                out<=15'b111100010100110;
            else if(A==8'd35)
                out<=15'b111011000011101;
            else if(A==8'd36)
                out<=15'b111110101010110;
            else if(A==8'd37)
                out<=15'b111101011001101;
            else if(A==8'd38)
                out<=15'b111100111001111;
            else if(A==8'd39)
                out<=15'b111011101000110;
            else if(A==8'd40)
                out<=15'b000000000101000;
            else if(A==8'd41)
                out<=15'b111110110011111;
            else if(A==8'd42)
                out<=15'b111110010100001;
            else if(A==8'd43)
                out<=15'b111101000011000;
            else if(A==8'd44)
                out<=15'b000000101010001;
            else if(A==8'd45)
                out<=15'b111111011001000;
            else if(A==8'd46)
                out<=15'b111110111001010;
            else if(A==8'd47)
                out<=15'b111101101000001;
            else if(A==8'd48)
                out<=15'b111110010010001;
            else if(A==8'd49)
                out<=15'b111101000001000;
            else if(A==8'd50)
                out<=15'b111100100001010;
            else if(A==8'd51)
                out<=15'b111011010000001;
            else if(A==8'd52)
                out<=15'b111110110111010;
            else if(A==8'd53)
                out<=15'b111101100110001;
            else if(A==8'd54)
                out<=15'b111101000110011;
            else if(A==8'd55)
                out<=15'b111011110101010;
            else if(A==8'd56)
                out<=15'b000000010001100;
            else if(A==8'd57)
                out<=15'b111111000000011;
            else if(A==8'd58)
                out<=15'b111110100000101;
            else if(A==8'd59)
                out<=15'b111101001111100;
            else if(A==8'd60)
                out<=15'b000000110110101;
            else if(A==8'd61)
                out<=15'b111111100101100;
            else if(A==8'd62)
                out<=15'b111111000101110;
            else if(A==8'd63)
                out<=15'b111101110100101;
            else if(A==8'd64)
                out<=15'b111111000011110;
            else if(A==8'd65)
                out<=15'b111101110010101;
            else if(A==8'd66)
                out<=15'b111101010010111;
            else if(A==8'd67)
                out<=15'b111100000001110;
            else if(A==8'd68)
                out<=15'b111111101000111;
            else if(A==8'd69)
                out<=15'b111110010111110;
            else if(A==8'd70)
                out<=15'b111101111000000;
            else if(A==8'd71)
                out<=15'b111100100110111;
            else if(A==8'd72)
                out<=15'b000001000011001;
            else if(A==8'd73)
                out<=15'b111111110010000;
            else if(A==8'd74)
                out<=15'b111111010010010;
            else if(A==8'd75)
                out<=15'b111110000001001;
            else if(A==8'd76)
                out<=15'b000001101000010;
            else if(A==8'd77)
                out<=15'b000000010111001;
            else if(A==8'd78)
                out<=15'b111111110111011;
            else if(A==8'd79)
                out<=15'b111110100110010;
            else if(A==8'd80)
                out<=15'b111111010000010;
            else if(A==8'd81)
                out<=15'b111101111111001;
            else if(A==8'd82)
                out<=15'b111101011111011;
            else if(A==8'd83)
                out<=15'b111100001110010;
            else if(A==8'd84)
                out<=15'b111111110101011;
            else if(A==8'd85)
                out<=15'b111110100100010;
            else if(A==8'd86)
                out<=15'b111110000100100;
            else if(A==8'd87)
                out<=15'b111100110011011;
            else if(A==8'd88)
                out<=15'b000001001111101;
            else if(A==8'd89)
                out<=15'b111111111110100;
            else if(A==8'd90)
                out<=15'b111111011110110;
            else if(A==8'd91)
                out<=15'b111110001101101;
            else if(A==8'd92)
                out<=15'b000001110100110;
            else if(A==8'd93)
                out<=15'b000000100011101;
            else if(A==8'd94)
                out<=15'b000000000011111;
            else if(A==8'd95)
                out<=15'b111110110010110;
            else if(A==8'd96)
                out<=15'b111101001001011;
            else if(A==8'd97)
                out<=15'b111011111000010;
            else if(A==8'd98)
                out<=15'b111011011000100;
            else if(A==8'd99)
                out<=15'b111010000111011;
            else if(A==8'd100)
                out<=15'b111101101110100;
            else if(A==8'd101)
                out<=15'b111100011101011;
            else if(A==8'd102)
                out<=15'b111011111101101;
            else if(A==8'd103)
                out<=15'b111010101100100;
            else if(A==8'd104)
                out<=15'b111111001000110;
            else if(A==8'd105)
                out<=15'b111101110111101;
            else if(A==8'd106)
                out<=15'b111101010111111;
            else if(A==8'd107)
                out<=15'b111100000110110;
            else if(A==8'd108)
                out<=15'b111111101101111;
            else if(A==8'd109)
                out<=15'b111110011100110;
            else if(A==8'd110)
                out<=15'b111101111101000;
            else if(A==8'd111)
                out<=15'b111100101011111;
            else if(A==8'd112)
                out<=15'b111101010101111;
            else if(A==8'd113)
                out<=15'b111100000100110;
            else if(A==8'd114)
                out<=15'b111011100101000;
            else if(A==8'd115)
                out<=15'b111010010011111;
            else if(A==8'd116)
                out<=15'b111101111011000;
            else if(A==8'd117)
                out<=15'b111100101001111;
            else if(A==8'd118)
                out<=15'b111100001010001;
            else if(A==8'd119)
                out<=15'b111010111001000;
            else if(A==8'd120)
                out<=15'b111111010101010;
            else if(A==8'd121)
                out<=15'b111110000100001;
            else if(A==8'd122)
                out<=15'b111101100100011;
            else if(A==8'd123)
                out<=15'b111100010011010;
            else if(A==8'd124)
                out<=15'b111111111010011;
            else if(A==8'd125)
                out<=15'b111110101001010;
            else if(A==8'd126)
                out<=15'b111110001001100;
            else if(A==8'd127)
                out<=15'b111100111000011;
            else if(A==8'd128)
                out<=15'b000001100010111;
            else if(A==8'd129)
                out<=15'b000000010001110;
            else if(A==8'd130)
                out<=15'b111111110010000;
            else if(A==8'd131)
                out<=15'b111110100000111;
            else if(A==8'd132)
                out<=15'b000010001000000;
            else if(A==8'd133)
                out<=15'b000000110110111;
            else if(A==8'd134)
                out<=15'b000000010111001;
            else if(A==8'd135)
                out<=15'b111111000110000;
            else if(A==8'd136)
                out<=15'b000011100010010;
            else if(A==8'd137)
                out<=15'b000010010001001;
            else if(A==8'd138)
                out<=15'b000001110001011;
            else if(A==8'd139)
                out<=15'b000000100000010;
            else if(A==8'd140)
                out<=15'b000100000111011;
            else if(A==8'd141)
                out<=15'b000010110110010;
            else if(A==8'd142)
                out<=15'b000010010110100;
            else if(A==8'd143)
                out<=15'b000001000101011;
            else if(A==8'd144)
                out<=15'b000001101111011;
            else if(A==8'd145)
                out<=15'b000000011110010;
            else if(A==8'd146)
                out<=15'b111111111110100;
            else if(A==8'd147)
                out<=15'b111110101101011;
            else if(A==8'd148)
                out<=15'b000010010100100;
            else if(A==8'd149)
                out<=15'b000001000011011;
            else if(A==8'd150)
                out<=15'b000000100011101;
            else if(A==8'd151)
                out<=15'b111111010010100;
            else if(A==8'd152)
                out<=15'b000011101110110;
            else if(A==8'd153)
                out<=15'b000010011101101;
            else if(A==8'd154)
                out<=15'b000001111101111;
            else if(A==8'd155)
                out<=15'b000000101100110;
            else if(A==8'd156)
                out<=15'b000100010011111;
            else if(A==8'd157)
                out<=15'b000011000010110;
            else if(A==8'd158)
                out<=15'b000010100011000;
            else if(A==8'd159)
                out<=15'b000001010001111;
            else if(A==8'd160)
                out<=15'b111111101000100;
            else if(A==8'd161)
                out<=15'b111110010111011;
            else if(A==8'd162)
                out<=15'b111101110111101;
            else if(A==8'd163)
                out<=15'b111100100110100;
            else if(A==8'd164)
                out<=15'b000000001101101;
            else if(A==8'd165)
                out<=15'b111110111100100;
            else if(A==8'd166)
                out<=15'b111110011100110;
            else if(A==8'd167)
                out<=15'b111101001011101;
            else if(A==8'd168)
                out<=15'b000001100111111;
            else if(A==8'd169)
                out<=15'b000000010110110;
            else if(A==8'd170)
                out<=15'b111111110111000;
            else if(A==8'd171)
                out<=15'b111110100101111;
            else if(A==8'd172)
                out<=15'b000010001101000;
            else if(A==8'd173)
                out<=15'b000000111011111;
            else if(A==8'd174)
                out<=15'b000000011100001;
            else if(A==8'd175)
                out<=15'b111111001011000;
            else if(A==8'd176)
                out<=15'b111111110101000;
            else if(A==8'd177)
                out<=15'b111110100011111;
            else if(A==8'd178)
                out<=15'b111110000100001;
            else if(A==8'd179)
                out<=15'b111100110011000;
            else if(A==8'd180)
                out<=15'b000000011010001;
            else if(A==8'd181)
                out<=15'b111111001001000;
            else if(A==8'd182)
                out<=15'b111110101001010;
            else if(A==8'd183)
                out<=15'b111101011000001;
            else if(A==8'd184)
                out<=15'b000001110100011;
            else if(A==8'd185)
                out<=15'b000000100011010;
            else if(A==8'd186)
                out<=15'b000000000011100;
            else if(A==8'd187)
                out<=15'b111110110010011;
            else if(A==8'd188)
                out<=15'b000010011001100;
            else if(A==8'd189)
                out<=15'b000001001000011;
            else if(A==8'd190)
                out<=15'b000000101000101;
            else if(A==8'd191)
                out<=15'b111111010111100;
            else if(A==8'd192)
                out<=15'b000000100110101;
            else if(A==8'd193)
                out<=15'b111111010101100;
            else if(A==8'd194)
                out<=15'b111110110101110;
            else if(A==8'd195)
                out<=15'b111101100100101;
            else if(A==8'd196)
                out<=15'b000001001011110;
            else if(A==8'd197)
                out<=15'b111111111010101;
            else if(A==8'd198)
                out<=15'b111111011010111;
            else if(A==8'd199)
                out<=15'b111110001001110;
            else if(A==8'd200)
                out<=15'b000010100110000;
            else if(A==8'd201)
                out<=15'b000001010100111;
            else if(A==8'd202)
                out<=15'b000000110101001;
            else if(A==8'd203)
                out<=15'b111111100100000;
            else if(A==8'd204)
                out<=15'b000011001011001;
            else if(A==8'd205)
                out<=15'b000001111010000;
            else if(A==8'd206)
                out<=15'b000001011010010;
            else if(A==8'd207)
                out<=15'b000000001001001;
            else if(A==8'd208)
                out<=15'b000000110011001;
            else if(A==8'd209)
                out<=15'b111111100010000;
            else if(A==8'd210)
                out<=15'b111111000010010;
            else if(A==8'd211)
                out<=15'b111101110001001;
            else if(A==8'd212)
                out<=15'b000001011000010;
            else if(A==8'd213)
                out<=15'b000000000111001;
            else if(A==8'd214)
                out<=15'b111111100111011;
            else if(A==8'd215)
                out<=15'b111110010110010;
            else if(A==8'd216)
                out<=15'b000010110010100;
            else if(A==8'd217)
                out<=15'b000001100001011;
            else if(A==8'd218)
                out<=15'b000001000001101;
            else if(A==8'd219)
                out<=15'b111111110000100;
            else if(A==8'd220)
                out<=15'b000011010111101;
            else if(A==8'd221)
                out<=15'b000010000110100;
            else if(A==8'd222)
                out<=15'b000001100110110;
            else if(A==8'd223)
                out<=15'b000000010101101;
            else if(A==8'd224)
                out<=15'b111110101100010;
            else if(A==8'd225)
                out<=15'b111101011011001;
            else if(A==8'd226)
                out<=15'b111100111011011;
            else if(A==8'd227)
                out<=15'b111011101010010;
            else if(A==8'd228)
                out<=15'b111111010001011;
            else if(A==8'd229)
                out<=15'b111110000000010;
            else if(A==8'd230)
                out<=15'b111101100000100;
            else if(A==8'd231)
                out<=15'b111100001111011;
            else if(A==8'd232)
                out<=15'b000000101011101;
            else if(A==8'd233)
                out<=15'b111111011010100;
            else if(A==8'd234)
                out<=15'b111110111010110;
            else if(A==8'd235)
                out<=15'b111101101001101;
            else if(A==8'd236)
                out<=15'b000001010000110;
            else if(A==8'd237)
                out<=15'b111111111111101;
            else if(A==8'd238)
                out<=15'b111111011111111;
            else if(A==8'd239)
                out<=15'b111110001110110;
            else if(A==8'd240)
                out<=15'b111110111000110;
            else if(A==8'd241)
                out<=15'b111101100111101;
            else if(A==8'd242)
                out<=15'b111101000111111;
            else if(A==8'd243)
                out<=15'b111011110110110;
            else if(A==8'd244)
                out<=15'b111111011101111;
            else if(A==8'd245)
                out<=15'b111110001100110;
            else if(A==8'd246)
                out<=15'b111101101101000;
            else if(A==8'd247)
                out<=15'b111100011011111;
            else if(A==8'd248)
                out<=15'b000000111000001;
            else if(A==8'd249)
                out<=15'b111111100111000;
            else if(A==8'd250)
                out<=15'b111111000111010;
            else if(A==8'd251)
                out<=15'b111101110110001;
            else if(A==8'd252)
                out<=15'b000001011101010;
            else if(A==8'd253)
                out<=15'b000000001100001;
            else if(A==8'd254)
                out<=15'b111111101100011;
            else
                out<=15'b111110011011010;      
        end
        
    else if(k==2)
        begin
            if(A==8'd0)
                out<=15'b000000000000000;
            else if(A==8'd1)
                out<=15'b111110001111001;
            else if(A==8'd2)
                out<=15'b000000001100100;
            else if(A==8'd3)
                out<=15'b111110011011101;
            else if(A==8'd4)
                out<=15'b000001100010111;
            else if(A==8'd5)
                out<=15'b111111110010000;
            else if(A==8'd6)
                out<=15'b000001101111011;
            else if(A==8'd7)
                out<=15'b111111111110100;
            else if(A==8'd8)
                out<=15'b111110000101101;
            else if(A==8'd9)
                out<=15'b111100010100110;
            else if(A==8'd10)
                out<=15'b111110010010001;
            else if(A==8'd11)
                out<=15'b111100100001010;
            else if(A==8'd12)
                out<=15'b111111101000100;
            else if(A==8'd13)
                out<=15'b111101110111101;
            else if(A==8'd14)
                out<=15'b111111110101000;
            else if(A==8'd15)
                out<=15'b111110000100001;
            else if(A==8'd16)
                out<=15'b000000100101001;
            else if(A==8'd17)
                out<=15'b111110110100010;
            else if(A==8'd18)
                out<=15'b000000110001101;
            else if(A==8'd19)
                out<=15'b111111000000110;
            else if(A==8'd20)
                out<=15'b000010001000000;
            else if(A==8'd21)
                out<=15'b000000010111001;
            else if(A==8'd22)
                out<=15'b000010010100100;
            else if(A==8'd23)
                out<=15'b000000100011101;
            else if(A==8'd24)
                out<=15'b111110101010110;
            else if(A==8'd25)
                out<=15'b111100111001111;
            else if(A==8'd26)
                out<=15'b111110110111010;
            else if(A==8'd27)
                out<=15'b111101000110011;
            else if(A==8'd28)
                out<=15'b000000001101101;
            else if(A==8'd29)
                out<=15'b111110011100110;
            else if(A==8'd30)
                out<=15'b000000011010001;
            else if(A==8'd31)
                out<=15'b111110101001010;
            else if(A==8'd32)
                out<=15'b000001010001001;
            else if(A==8'd33)
                out<=15'b111111100000010;
            else if(A==8'd34)
                out<=15'b000001011101101;
            else if(A==8'd35)
                out<=15'b111111101100110;
            else if(A==8'd36)
                out<=15'b000010110100000;
            else if(A==8'd37)
                out<=15'b000001000011001;
            else if(A==8'd38)
                out<=15'b000011000000100;
            else if(A==8'd39)
                out<=15'b000001001111101;
            else if(A==8'd40)
                out<=15'b111111010110110;
            else if(A==8'd41)
                out<=15'b111101100101111;
            else if(A==8'd42)
                out<=15'b111111100011010;
            else if(A==8'd43)
                out<=15'b111101110010011;
            else if(A==8'd44)
                out<=15'b000000111001101;
            else if(A==8'd45)
                out<=15'b111111001000110;
            else if(A==8'd46)
                out<=15'b000001000110001;
            else if(A==8'd47)
                out<=15'b111111010101010;
            else if(A==8'd48)
                out<=15'b000001110110010;
            else if(A==8'd49)
                out<=15'b000000000101011;
            else if(A==8'd50)
                out<=15'b000010000010110;
            else if(A==8'd51)
                out<=15'b000000010001111;
            else if(A==8'd52)
                out<=15'b000011011001001;
            else if(A==8'd53)
                out<=15'b000001101000010;
            else if(A==8'd54)
                out<=15'b000011100101101;
            else if(A==8'd55)
                out<=15'b000001110100110;
            else if(A==8'd56)
                out<=15'b111111111011111;
            else if(A==8'd57)
                out<=15'b111110001011000;
            else if(A==8'd58)
                out<=15'b000000001000011;
            else if(A==8'd59)
                out<=15'b111110010111100;
            else if(A==8'd60)
                out<=15'b000001011110110;
            else if(A==8'd61)
                out<=15'b111111101101111;
            else if(A==8'd62)
                out<=15'b000001101011010;
            else if(A==8'd63)
                out<=15'b111111111010011;
            else if(A==8'd64)
                out<=15'b111110000000101;
            else if(A==8'd65)
                out<=15'b111100001111110;
            else if(A==8'd66)
                out<=15'b111110001101001;
            else if(A==8'd67)
                out<=15'b111100011100010;
            else if(A==8'd68)
                out<=15'b111111100011100;
            else if(A==8'd69)
                out<=15'b111101110010101;
            else if(A==8'd70)
                out<=15'b111111110000000;
            else if(A==8'd71)
                out<=15'b111101111111001;
            else if(A==8'd72)
                out<=15'b111100000110010;
            else if(A==8'd73)
                out<=15'b111010010101011;
            else if(A==8'd74)
                out<=15'b111100010010110;
            else if(A==8'd75)
                out<=15'b111010100001111;
            else if(A==8'd76)
                out<=15'b111101101001001;
            else if(A==8'd77)
                out<=15'b111011111000010;
            else if(A==8'd78)
                out<=15'b111101110101101;
            else if(A==8'd79)
                out<=15'b111100000100110;
            else if(A==8'd80)
                out<=15'b111110100101110;
            else if(A==8'd81)
                out<=15'b111100110100111;
            else if(A==8'd82)
                out<=15'b111110110010010;
            else if(A==8'd83)
                out<=15'b111101000001011;
            else if(A==8'd84)
                out<=15'b000000001000101;
            else if(A==8'd85)
                out<=15'b111110010111110;
            else if(A==8'd86)
                out<=15'b000000010101001;
            else if(A==8'd87)
                out<=15'b111110100100010;
            else if(A==8'd88)
                out<=15'b111100101011011;
            else if(A==8'd89)
                out<=15'b111010111010100;
            else if(A==8'd90)
                out<=15'b111100110111111;
            else if(A==8'd91)
                out<=15'b111011000111000;
            else if(A==8'd92)
                out<=15'b111110001110010;
            else if(A==8'd93)
                out<=15'b111100011101011;
            else if(A==8'd94)
                out<=15'b111110011010110;
            else if(A==8'd95)
                out<=15'b111100101001111;
            else if(A==8'd96)
                out<=15'b111111010001110;
            else if(A==8'd97)
                out<=15'b111101100000111;
            else if(A==8'd98)
                out<=15'b111111011110010;
            else if(A==8'd99)
                out<=15'b111101101101011;
            else if(A==8'd100)
                out<=15'b000000110100101;
            else if(A==8'd101)
                out<=15'b111111000011110;
            else if(A==8'd102)
                out<=15'b000001000001001;
            else if(A==8'd103)
                out<=15'b111111010000010;
            else if(A==8'd104)
                out<=15'b111101010111011;
            else if(A==8'd105)
                out<=15'b111011100110100;
            else if(A==8'd106)
                out<=15'b111101100011111;
            else if(A==8'd107)
                out<=15'b111011110011000;
            else if(A==8'd108)
                out<=15'b111110111010010;
            else if(A==8'd109)
                out<=15'b111101001001011;
            else if(A==8'd110)
                out<=15'b111111000110110;
            else if(A==8'd111)
                out<=15'b111101010101111;
            else if(A==8'd112)
                out<=15'b111111110110111;
            else if(A==8'd113)
                out<=15'b111110000110000;
            else if(A==8'd114)
                out<=15'b000000000011011;
            else if(A==8'd115)
                out<=15'b111110010010100;
            else if(A==8'd116)
                out<=15'b000001011001110;
            else if(A==8'd117)
                out<=15'b111111101000111;
            else if(A==8'd118)
                out<=15'b000001100110010;
            else if(A==8'd119)
                out<=15'b111111110101011;
            else if(A==8'd120)
                out<=15'b111101111100100;
            else if(A==8'd121)
                out<=15'b111100001011101;
            else if(A==8'd122)
                out<=15'b111110001001000;
            else if(A==8'd123)
                out<=15'b111100011000001;
            else if(A==8'd124)
                out<=15'b111111011111011;
            else if(A==8'd125)
                out<=15'b111101101110100;
            else if(A==8'd126)
                out<=15'b111111101011111;
            else if(A==8'd127)
                out<=15'b111101111011000;
            else if(A==8'd128)
                out<=15'b000000111100010;
            else if(A==8'd129)
                out<=15'b111111001011011;
            else if(A==8'd130)
                out<=15'b000001001000110;
            else if(A==8'd131)
                out<=15'b111111010111111;
            else if(A==8'd132)
                out<=15'b000010011111001;
            else if(A==8'd133)
                out<=15'b000000101110010;
            else if(A==8'd134)
                out<=15'b000010101011101;
            else if(A==8'd135)
                out<=15'b000000111010110;
            else if(A==8'd136)
                out<=15'b111111000001111;
            else if(A==8'd137)
                out<=15'b111101010001000;
            else if(A==8'd138)
                out<=15'b111111001110011;
            else if(A==8'd139)
                out<=15'b111101011101100;
            else if(A==8'd140)
                out<=15'b000000100100110;
            else if(A==8'd141)
                out<=15'b111110110011111;
            else if(A==8'd142)
                out<=15'b000000110001010;
            else if(A==8'd143)
                out<=15'b111111000000011;
            else if(A==8'd144)
                out<=15'b000001100001011;
            else if(A==8'd145)
                out<=15'b111111110000100;
            else if(A==8'd146)
                out<=15'b000001101101111;
            else if(A==8'd147)
                out<=15'b111111111101000;
            else if(A==8'd148)
                out<=15'b000011000100010;
            else if(A==8'd149)
                out<=15'b000001010011011;
            else if(A==8'd150)
                out<=15'b000011010000110;
            else if(A==8'd151)
                out<=15'b000001011111111;
            else if(A==8'd152)
                out<=15'b111111100111000;
            else if(A==8'd153)
                out<=15'b111101110110001;
            else if(A==8'd154)
                out<=15'b111111110011100;
            else if(A==8'd155)
                out<=15'b111110000010101;
            else if(A==8'd156)
                out<=15'b000001001001111;
            else if(A==8'd157)
                out<=15'b111111011001000;
            else if(A==8'd158)
                out<=15'b000001010110011;
            else if(A==8'd159)
                out<=15'b111111100101100;
            else if(A==8'd160)
                out<=15'b000010001101011;
            else if(A==8'd161)
                out<=15'b000000011100100;
            else if(A==8'd162)
                out<=15'b000010011001111;
            else if(A==8'd163)
                out<=15'b000000101001000;
            else if(A==8'd164)
                out<=15'b000011110000010;
            else if(A==8'd165)
                out<=15'b000001111111011;
            else if(A==8'd166)
                out<=15'b000011111100110;
            else if(A==8'd167)
                out<=15'b000010001011111;
            else if(A==8'd168)
                out<=15'b000000010011000;
            else if(A==8'd169)
                out<=15'b111110100010001;
            else if(A==8'd170)
                out<=15'b000000011111100;
            else if(A==8'd171)
                out<=15'b111110101110101;
            else if(A==8'd172)
                out<=15'b000001110101111;
            else if(A==8'd173)
                out<=15'b000000000101000;
            else if(A==8'd174)
                out<=15'b000010000010011;
            else if(A==8'd175)
                out<=15'b000000010001100;
            else if(A==8'd176)
                out<=15'b000010110010100;
            else if(A==8'd177)
                out<=15'b000001000001101;
            else if(A==8'd178)
                out<=15'b000010111111000;
            else if(A==8'd179)
                out<=15'b000001001110001;
            else if(A==8'd180)
                out<=15'b000100010101011;
            else if(A==8'd181)
                out<=15'b000010100100100;
            else if(A==8'd182)
                out<=15'b000100100001111;
            else if(A==8'd183)
                out<=15'b000010110001000;
            else if(A==8'd184)
                out<=15'b000000111000001;
            else if(A==8'd185)
                out<=15'b111111000111010;
            else if(A==8'd186)
                out<=15'b000001000100101;
            else if(A==8'd187)
                out<=15'b111111010011110;
            else if(A==8'd188)
                out<=15'b000010011011000;
            else if(A==8'd189)
                out<=15'b000000101010001;
            else if(A==8'd190)
                out<=15'b000010100111100;
            else if(A==8'd191)
                out<=15'b000000110110101;
            else if(A==8'd192)
                out<=15'b111110111100111;
            else if(A==8'd193)
                out<=15'b111101001100000;
            else if(A==8'd194)
                out<=15'b111111001001011;
            else if(A==8'd195)
                out<=15'b111101011000100;
            else if(A==8'd196)
                out<=15'b000000011111110;
            else if(A==8'd197)
                out<=15'b111110101110111;
            else if(A==8'd198)
                out<=15'b000000101100010;
            else if(A==8'd199)
                out<=15'b111110111011011;
            else if(A==8'd200)
                out<=15'b111101000010100;
            else if(A==8'd201)
                out<=15'b111011010001101;
            else if(A==8'd202)
                out<=15'b111101001111000;
            else if(A==8'd203)
                out<=15'b111011011110001;
            else if(A==8'd204)
                out<=15'b111110100101011;
            else if(A==8'd205)
                out<=15'b111100110100100;
            else if(A==8'd206)
                out<=15'b111110110001111;
            else if(A==8'd207)
                out<=15'b111101000001000;
            else if(A==8'd208)
                out<=15'b111111100010000;
            else if(A==8'd209)
                out<=15'b111101110001001;
            else if(A==8'd210)
                out<=15'b111111101110100;
            else if(A==8'd211)
                out<=15'b111101111101101;
            else if(A==8'd212)
                out<=15'b000001000100111;
            else if(A==8'd213)
                out<=15'b111111010100000;
            else if(A==8'd214)
                out<=15'b000001010001011;
            else if(A==8'd215)
                out<=15'b111111100000100;
            else if(A==8'd216)
                out<=15'b111101100111101;
            else if(A==8'd217)
                out<=15'b111011110110110;
            else if(A==8'd218)
                out<=15'b111101110100001;
            else if(A==8'd219)
                out<=15'b111100000011010;
            else if(A==8'd220)
                out<=15'b111111001010100;
            else if(A==8'd221)
                out<=15'b111101011001101;
            else if(A==8'd222)
                out<=15'b111111010111000;
            else if(A==8'd223)
                out<=15'b111101100110001;
            else if(A==8'd224)
                out<=15'b000000001110000;
            else if(A==8'd225)
                out<=15'b111110011101001;
            else if(A==8'd226)
                out<=15'b000000011010100;
            else if(A==8'd227)
                out<=15'b111110101001101;
            else if(A==8'd228)
                out<=15'b000001110000111;
            else if(A==8'd229)
                out<=15'b000000000000000;
            else if(A==8'd230)
                out<=15'b000001111101011;
            else if(A==8'd231)
                out<=15'b000000001100100;
            else if(A==8'd232)
                out<=15'b111110010011101;
            else if(A==8'd233)
                out<=15'b111100100010110;
            else if(A==8'd234)
                out<=15'b111110100000001;
            else if(A==8'd235)
                out<=15'b111100101111010;
            else if(A==8'd236)
                out<=15'b111111110110100;
            else if(A==8'd237)
                out<=15'b111110000101101;
            else if(A==8'd238)
                out<=15'b000000000011000;
            else if(A==8'd239)
                out<=15'b111110010010001;
            else if(A==8'd240)
                out<=15'b000000110011001;
            else if(A==8'd241)
                out<=15'b111111000010010;
            else if(A==8'd242)
                out<=15'b000000111111101;
            else if(A==8'd243)
                out<=15'b111111001110110;
            else if(A==8'd244)
                out<=15'b000010010110000;
            else if(A==8'd245)
                out<=15'b000000100101001;
            else if(A==8'd246)
                out<=15'b000010100010100;
            else if(A==8'd247)
                out<=15'b000000110001101;
            else if(A==8'd248)
                out<=15'b111110111000110;
            else if(A==8'd249)
                out<=15'b111101000111111;
            else if(A==8'd250)
                out<=15'b111111000101010;
            else if(A==8'd251)
                out<=15'b111101010100011;
            else if(A==8'd252)
                out<=15'b000000011011101;
            else if(A==8'd253)
                out<=15'b111110101010110;
            else if(A==8'd254)
                out<=15'b000000101000001;
            else 
                out<=15'b111110110111010;             
        end
        
     //else if(k==3)
     else 
        begin
            if(A==8'd0)
                out<=15'b000000000000000;
            else if(A==8'd1)
                out<=15'b111110000000101;
            else if(A==8'd2)
                out<=15'b000001111010011;
            else if(A==8'd3)
                out<=15'b111111111011000;
            else if(A==8'd4)
                out<=15'b111110001111001;
            else if(A==8'd5)
                out<=15'b111100001111110;
            else if(A==8'd6)
                out<=15'b000000001001100;
            else if(A==8'd7)
                out<=15'b111110001010001;
            else if(A==8'd8)
                out<=15'b000001100010111;
            else if(A==8'd9)
                out<=15'b111111100011100;
            else if(A==8'd10)
                out<=15'b000011011101010;
            else if(A==8'd11)
                out<=15'b000001011101111;
            else if(A==8'd12)
                out<=15'b111111110010000;
            else if(A==8'd13)
                out<=15'b111101110010101;
            else if(A==8'd14)
                out<=15'b000001101100011;
            else if(A==8'd15)
                out<=15'b111111101101000;
            else if(A==8'd16)
                out<=15'b111110101110111;
            else if(A==8'd17)
                out<=15'b111100101111100;
            else if(A==8'd18)
                out<=15'b000000101001010;
            else if(A==8'd19)
                out<=15'b111110101001111;
            else if(A==8'd20)
                out<=15'b111100111110000;
            else if(A==8'd21)
                out<=15'b111010111110101;
            else if(A==8'd22)
                out<=15'b111110111000011;
            else if(A==8'd23)
                out<=15'b111100111001000;
            else if(A==8'd24)
                out<=15'b000000010001110;
            else if(A==8'd25)
                out<=15'b111110010010011;
            else if(A==8'd26)
                out<=15'b000010001100001;
            else if(A==8'd27)
                out<=15'b000000001100110;
            else if(A==8'd28)
                out<=15'b111110100000111;
            else if(A==8'd29)
                out<=15'b111100100001100;
            else if(A==8'd30)
                out<=15'b000000011011010;
            else if(A==8'd31)
                out<=15'b111110011011111;
            else if(A==8'd32)
                out<=15'b000000111100010;
            else if(A==8'd33)
                out<=15'b111110111100111;
            else if(A==8'd34)
                out<=15'b000010110110101;
            else if(A==8'd35)
                out<=15'b000000110111010;
            else if(A==8'd36)
                out<=15'b111111001011011;
            else if(A==8'd37)
                out<=15'b111101001100000;
            else if(A==8'd38)
                out<=15'b000001000101110;
            else if(A==8'd39)
                out<=15'b111111000110011;
            else if(A==8'd40)
                out<=15'b000010011111001;
            else if(A==8'd41)
                out<=15'b000000011111110;
            else if(A==8'd42)
                out<=15'b000100011001100;
            else if(A==8'd43)
                out<=15'b000010011010001;
            else if(A==8'd44)
                out<=15'b000000101110010;
            else if(A==8'd45)
                out<=15'b111110101110111;
            else if(A==8'd46)
                out<=15'b000010101000101;
            else if(A==8'd47)
                out<=15'b000000101001010;
            else if(A==8'd48)
                out<=15'b111111101011001;
            else if(A==8'd49)
                out<=15'b111101101011110;
            else if(A==8'd50)
                out<=15'b000001100101100;
            else if(A==8'd51)
                out<=15'b111111100110001;
            else if(A==8'd52)
                out<=15'b111101111010010;
            else if(A==8'd53)
                out<=15'b111011111010111;
            else if(A==8'd54)
                out<=15'b111111110100101;
            else if(A==8'd55)
                out<=15'b111101110101010;
            else if(A==8'd56)
                out<=15'b000001001110000;
            else if(A==8'd57)
                out<=15'b111111001110101;
            else if(A==8'd58)
                out<=15'b000011001000011;
            else if(A==8'd59)
                out<=15'b000001001001000;
            else if(A==8'd60)
                out<=15'b111111011101001;
            else if(A==8'd61)
                out<=15'b111101011101110;
            else if(A==8'd62)
                out<=15'b000001010111100;
            else if(A==8'd63)
                out<=15'b111111011000001;
            else if(A==8'd64)
                out<=15'b111111011010111;
            else if(A==8'd65)
                out<=15'b111101011011100;
            else if(A==8'd66)
                out<=15'b000001010101010;
            else if(A==8'd67)
                out<=15'b111111010101111;
            else if(A==8'd68)
                out<=15'b111101101010000;
            else if(A==8'd69)
                out<=15'b111011101010101;
            else if(A==8'd70)
                out<=15'b111111100100011;
            else if(A==8'd71)
                out<=15'b111101100101000;
            else if(A==8'd72)
                out<=15'b000000111101110;
            else if(A==8'd73)
                out<=15'b111110111110011;
            else if(A==8'd74)
                out<=15'b000010111000001;
            else if(A==8'd75)
                out<=15'b000000111000110;
            else if(A==8'd76)
                out<=15'b111111001100111;
            else if(A==8'd77)
                out<=15'b111101001101100;
            else if(A==8'd78)
                out<=15'b000001000111010;
            else if(A==8'd79)
                out<=15'b111111000111111;
            else if(A==8'd80)
                out<=15'b111110001001110;
            else if(A==8'd81)
                out<=15'b111100001010011;
            else if(A==8'd82)
                out<=15'b000000000100001;
            else if(A==8'd83)
                out<=15'b111110000100110;
            else if(A==8'd84)
                out<=15'b111100011000111;
            else if(A==8'd85)
                out<=15'b111010011001100;
            else if(A==8'd86)
                out<=15'b111110010011010;
            else if(A==8'd87)
                out<=15'b111100010011111;
            else if(A==8'd88)
                out<=15'b111111101100101;
            else if(A==8'd89)
                out<=15'b111101101101010;
            else if(A==8'd90)
                out<=15'b000001100111000;
            else if(A==8'd91)
                out<=15'b111111100111101;
            else if(A==8'd92)
                out<=15'b111101111011110;
            else if(A==8'd93)
                out<=15'b111011111100011;
            else if(A==8'd94)
                out<=15'b111111110110001;
            else if(A==8'd95)
                out<=15'b111101110110110;
            else if(A==8'd96)
                out<=15'b000000010111001;
            else if(A==8'd97)
                out<=15'b111110010111110;
            else if(A==8'd98)
                out<=15'b000010010001100;
            else if(A==8'd99)
                out<=15'b000000010010001;
            else if(A==8'd100)
                out<=15'b111110100110010;
            else if(A==8'd101)
                out<=15'b111100100110111;
            else if(A==8'd102)
                out<=15'b000000100000101;
            else if(A==8'd103)
                out<=15'b111110100001010;
            else if(A==8'd104)
                out<=15'b000001111010000;
            else if(A==8'd105)
                out<=15'b111111111010101;
            else if(A==8'd106)
                out<=15'b000011110100011;
            else if(A==8'd107)
                out<=15'b000001110101000;
            else if(A==8'd108)
                out<=15'b000000001001001;
            else if(A==8'd109)
                out<=15'b111110001001110;
            else if(A==8'd110)
                out<=15'b000010000011100;
            else if(A==8'd111)
                out<=15'b000000000100001;
            else if(A==8'd112)
                out<=15'b111111000110000;
            else if(A==8'd113)
                out<=15'b111101000110101;
            else if(A==8'd114)
                out<=15'b000001000000011;
            else if(A==8'd115)
                out<=15'b111111000001000;
            else if(A==8'd116)
                out<=15'b111101010101001;
            else if(A==8'd117)
                out<=15'b111011010101110;
            else if(A==8'd118)
                out<=15'b111111001111100;
            else if(A==8'd119)
                out<=15'b111101010000001;
            else if(A==8'd120)
                out<=15'b000000101000111;
            else if(A==8'd121)
                out<=15'b111110101001100;
            else if(A==8'd122)
                out<=15'b000010100011010;
            else if(A==8'd123)
                out<=15'b000000100011111;
            else if(A==8'd124)
                out<=15'b111110111000000;
            else if(A==8'd125)
                out<=15'b111100111000101;
            else if(A==8'd126)
                out<=15'b000000110010011;
            else if(A==8'd127)
                out<=15'b111110110011000;
            else if(A==8'd128)
                out<=15'b000000001100100;
            else if(A==8'd129)
                out<=15'b111110001101001;
            else if(A==8'd130)
                out<=15'b000010000110111;
            else if(A==8'd131)
                out<=15'b000000000111100;
            else if(A==8'd132)
                out<=15'b111110011011101;
            else if(A==8'd133)
                out<=15'b111100011100010;
            else if(A==8'd134)
                out<=15'b000000010110000;
            else if(A==8'd135)
                out<=15'b111110010110101;
            else if(A==8'd136)
                out<=15'b000001101111011;
            else if(A==8'd137)
                out<=15'b111111110000000;
            else if(A==8'd138)
                out<=15'b000011101001110;
            else if(A==8'd139)
                out<=15'b000001101010011;
            else if(A==8'd140)
                out<=15'b111111111110100;
            else if(A==8'd141)
                out<=15'b111101111111001;
            else if(A==8'd142)
                out<=15'b000001111000111;
            else if(A==8'd143)
                out<=15'b111111111001100;
            else if(A==8'd144)
                out<=15'b111110111011011;
            else if(A==8'd145)
                out<=15'b111100111100000;
            else if(A==8'd146)
                out<=15'b000000110101110;
            else if(A==8'd147)
                out<=15'b111110110110011;
            else if(A==8'd148)
                out<=15'b111101001010100;
            else if(A==8'd149)
                out<=15'b111011001011001;
            else if(A==8'd150)
                out<=15'b111111000100111;
            else if(A==8'd151)
                out<=15'b111101000101100;
            else if(A==8'd152)
                out<=15'b000000011110010;
            else if(A==8'd153)
                out<=15'b111110011110111;
            else if(A==8'd154)
                out<=15'b000010011000101;
            else if(A==8'd155)
                out<=15'b000000011001010;
            else if(A==8'd156)
                out<=15'b111110101101011;
            else if(A==8'd157)
                out<=15'b111100101110000;
            else if(A==8'd158)
                out<=15'b000000100111110;
            else if(A==8'd159)
                out<=15'b111110101000011;
            else if(A==8'd160)
                out<=15'b000001001000110;
            else if(A==8'd161)
                out<=15'b111111001001011;
            else if(A==8'd162)
                out<=15'b000011000011001;
            else if(A==8'd163)
                out<=15'b000001000011110;
            else if(A==8'd164)
                out<=15'b111111010111111;
            else if(A==8'd165)
                out<=15'b111101011000100;
            else if(A==8'd166)
                out<=15'b000001010010010;
            else if(A==8'd167)
                out<=15'b111111010010111;
            else if(A==8'd168)
                out<=15'b000010101011101;
            else if(A==8'd169)
                out<=15'b000000101100010;
            else if(A==8'd170)
                out<=15'b000100100110000;
            else if(A==8'd171)
                out<=15'b000010100110101;
            else if(A==8'd172)
                out<=15'b000000111010110;
            else if(A==8'd173)
                out<=15'b111110111011011;
            else if(A==8'd174)
                out<=15'b000010110101001;
            else if(A==8'd175)
                out<=15'b000000110101110;
            else if(A==8'd176)
                out<=15'b111111110111101;
            else if(A==8'd177)
                out<=15'b111101111000010;
            else if(A==8'd178)
                out<=15'b000001110010000;
            else if(A==8'd179)
                out<=15'b111111110010101;
            else if(A==8'd180)
                out<=15'b111110000110110;
            else if(A==8'd181)
                out<=15'b111100000111011;
            else if(A==8'd182)
                out<=15'b000000000001001;
            else if(A==8'd183)
                out<=15'b111110000001110;
            else if(A==8'd184)
                out<=15'b000001011010100;
            else if(A==8'd185)
                out<=15'b111111011011001;
            else if(A==8'd186)
                out<=15'b000011010100111;
            else if(A==8'd187)
                out<=15'b000001010101100;
            else if(A==8'd188)
                out<=15'b111111101001101;
            else if(A==8'd189)
                out<=15'b111101101010010;
            else if(A==8'd190)
                out<=15'b000001100100000;
            else if(A==8'd191)
                out<=15'b111111100100101;
            else if(A==8'd192)
                out<=15'b111111100111011;
            else if(A==8'd193)
                out<=15'b111101101000000;
            else if(A==8'd194)
                out<=15'b000001100001110;
            else if(A==8'd195)
                out<=15'b111111100010011;
            else if(A==8'd196)
                out<=15'b111101110110100;
            else if(A==8'd197)
                out<=15'b111011110111001;
            else if(A==8'd198)
                out<=15'b111111110000111;
            else if(A==8'd199)
                out<=15'b111101110001100;
            else if(A==8'd200)
                out<=15'b000001001010010;
            else if(A==8'd201)
                out<=15'b111111001010111;
            else if(A==8'd202)
                out<=15'b000011000100101;
            else if(A==8'd203)
                out<=15'b000001000101010;
            else if(A==8'd204)
                out<=15'b111111011001011;
            else if(A==8'd205)
                out<=15'b111101011010000;
            else if(A==8'd206)
                out<=15'b000001010011110;
            else if(A==8'd207)
                out<=15'b111111010100011;
            else if(A==8'd208)
                out<=15'b111110010110010;
            else if(A==8'd209)
                out<=15'b111100010110111;
            else if(A==8'd210)
                out<=15'b000000010000101;
            else if(A==8'd211)
                out<=15'b111110010001010;
            else if(A==8'd212)
                out<=15'b111100100101011;
            else if(A==8'd213)
                out<=15'b111010100110000;
            else if(A==8'd214)
                out<=15'b111110011111110;
            else if(A==8'd215)
                out<=15'b111100100000011;
            else if(A==8'd216)
                out<=15'b111111111001001;
            else if(A==8'd217)
                out<=15'b111101111001110;
            else if(A==8'd218)
                out<=15'b000001110011100;
            else if(A==8'd219)
                out<=15'b111111110100001;
            else if(A==8'd220)
                out<=15'b111110001000010;
            else if(A==8'd221)
                out<=15'b111100001000111;
            else if(A==8'd222)
                out<=15'b000000000010101;
            else if(A==8'd223)
                out<=15'b111110000011010;
            else if(A==8'd224)
                out<=15'b000000100011101;
            else if(A==8'd225)
                out<=15'b111110100100010;
            else if(A==8'd226)
                out<=15'b000010011110000;
            else if(A==8'd227)
                out<=15'b000000011110101;
            else if(A==8'd228)
                out<=15'b111110110010110;
            else if(A==8'd229)
                out<=15'b111100110011011;
            else if(A==8'd230)
                out<=15'b000000101101001;
            else if(A==8'd231)
                out<=15'b111110101101110;
            else if(A==8'd232)
                out<=15'b000010000110100;
            else if(A==8'd233)
                out<=15'b000000000111001;
            else if(A==8'd234)
                out<=15'b000100000000111;
            else if(A==8'd235)
                out<=15'b000010000001100;
            else if(A==8'd236)
                out<=15'b000000010101101;
            else if(A==8'd237)
                out<=15'b111110010110010;
            else if(A==8'd238)
                out<=15'b000010010000000;
            else if(A==8'd239)
                out<=15'b000000010000101;
            else if(A==8'd240)
                out<=15'b111111010010100;
            else if(A==8'd241)
                out<=15'b111101010011001;
            else if(A==8'd242)
                out<=15'b000001001100111;
            else if(A==8'd243)
                out<=15'b111111001101100;
            else if(A==8'd244)
                out<=15'b111101100001101;
            else if(A==8'd245)
                out<=15'b111011100010010;
            else if(A==8'd246)
                out<=15'b111111011100000;
            else if(A==8'd247)
                out<=15'b111101011100101;
            else if(A==8'd248)
                out<=15'b000000110101011;
            else if(A==8'd249)
                out<=15'b111110110110000;
            else if(A==8'd250)
                out<=15'b000010101111110;
            else if(A==8'd251)
                out<=15'b000000110000011;
            else if(A==8'd252)
                out<=15'b111111000100100;
            else if(A==8'd253)
                out<=15'b111101000101001;
            else if(A==8'd254)
                out<=15'b000000111110111;
            else
                out<=15'b111110111111100;     
        end
       
             
end 
endmodule
